shifter_inst : shifter PORT MAP (
		data	 => data_sig,
		direction	 => direction_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
